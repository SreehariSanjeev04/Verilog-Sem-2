module main_circuit_tb;
parameter PRICE_1 = 4'b0001;
parameter PRICE_2 = 4'b0010;
parameter WEIGHT_THRESHOLD = 4'b0100;
parameter FAST_CHARGE_PRICE = 4'b0010;
parameter CHARGE_PRICE = 4'b0001;
parameter CHARGE_THRESHOLD = 4'b0100;
parameter HIGH_CAPACITY_PRICE = 4'b0010;
parameter SMALL_CAPACITY_PRICE = 4'b0001;
parameter CAPACITY_THRESHOLD = 4'b0100;
parameter PASSWORD = 4'b1101;
parameter WEIGHT = 4'b0110;
parameter PARK_SEQUENCE = 8'b11001100;
reg [3:0]user_password;
reg [7:0]additional;
reg [2:0]code;
reg [3:0]hours;
reg [3:0] temp;
reg [7:0] firePosition;
reg [3:0] duration;
reg [3:0] power;
reg [7:0] cash;
reg [3:0] capacity;
reg [3:0] card_number;
reg reverse;
wire password_matched,isPaidCash,isPaidCard;
wire [7:0] result,alarm_status;
main_circuit m1(PRICE_1,PRICE_2,WEIGHT_THRESHOLD,FAST_CHARGE_PRICE,CHARGE_PRICE,CHARGE_THRESHOLD,HIGH_CAPACITY_PRICE,SMALL_CAPACITY_PRICE,CAPACITY_THRESHOLD,temp,firePosition,duration,power,capacity,PASSWORD,user_password,WEIGHT,cash,card_number,PARK_SEQUENCE,additional,code,hours,reverse,password_matched,isPaidCash,isPaidCard,result,alarm_status);
initial begin
$monitor("CODE: %b\nPASSWORD MATCH:%b\nALARM STATUS: %b\nisPaidCash: %b\nisPaidCard: %b\nOutput: %b\n",code,password_matched,alarm_status,isPaidCash,isPaidCard,result);
user_password=4'b1100;
additional=8'b00100000;
code=3'b010;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0110;
cash=8'b10000000;
#10
user_password=4'b1100;
additional=8'b00100000;
code=3'b010;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b01000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0110;
cash=8'b00000000;
#10
user_password=4'b1101;
additional=8'b00000000;
code=3'b000;
temp=4'b0001;
hours=4'b0000;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0000;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0000;
cash=8'b00000000;
#10
user_password=4'b1101;
additional=8'b00100000;
code=3'b001;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0110;
cash=8'b00000000;
#10
user_password=4'b1101;
additional=8'b00100000;
code=3'b010;
temp=4'b0001;
hours=4'b0000;
firePosition=8'b00000000;
duration=4'b0000;
power=4'b0000;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0000;
cash=8'b00000000;
#10
user_password=4'b1101;
additional=8'b00100000;
code=3'b011;
temp=4'b0001;
hours=4'b0000;
firePosition=8'b00000000;
duration=4'b0000;
power=4'b0000;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0000;
cash=8'b10000000;
#10
user_password=4'b1101;
additional=8'b00100000;
code=3'b100;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0110;
cash=8'b10000000;
#10
user_password=4'b1101;
additional=8'b00100000;
code=3'b101;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0110;
cash=8'b10000000;
#10
user_password=4'b1101;
additional=8'b00000000;
code=3'b110;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0000;
cash=8'b00000000;
#10
user_password=4'b1101;
additional=8'b00100000;
code=3'b111;
temp=4'b0001;
hours=4'b0011;
firePosition=8'b00000000;
duration=4'b0101;
power=4'b0011;
capacity=4'b0000;
reverse=1'b0;
card_number=4'b0110;
cash=8'b10000000;

end
endmodule
